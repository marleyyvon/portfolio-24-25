module IM(Address, OUT);
input [31:0]Address;
output [31:0]OUT;
reg [31:0]data[255:0];
integer i;
initial begin
    // (1) Fill everything with NOPs
    for (i = 0; i < 256; i = i + 1) begin
      data[i] = 32'b0000_000000_000000_000000_0000000000;  // opcode=0000 = NOP
    end
    /*
    // LD   x5,  x10       // x5 ? M[x10]
    data[0]  = 32'b1110_000101_001010_000000_0000000000;

    // SVPC x6, 3          // x6 ? PC + 2  (loop start)
    data[1]  = 32'b1111_000110_0000000000000000000011;

    // SVPC x7, 12          // x7 ? PC + 7  (update "poop")
    data[2]  = 32'b1111_000111_0000000000000000001100;

    // INC  x11, x11, -1   // x11 ? x11 - 1 (loop counter--)
    data[3]  = 32'b0101_001011_001011_1111111111111111;
    data[4]  = 32'b0101_001011_001011_1111111111111111;
    // INC  x10, x10, 1    // x10 ? x10 + 1 (pointer++)
    data[5] = 32'b0101_001010_001010_0000000000000001;

    // LD   x28, x10       // x28 ? M[x10]
    data[6]  = 32'b1110_011100_001010_000000_0000000000;

    // SUB  x29, x5, x28   // x29 ? x5 - x28
    data[9]  = 32'b0111_011101_000101_011100_0000000000;

    // BRN  x7             // if N=1 (a[i]<poop) jump to update
    data[10]  = 32'b1011_000000_000111_000000_0000000000;

    // ADD  x5, x0, x28    // poop ? a[i]
    data[13]  = 32'b0100_000101_000000_011100_0000000000;

    // SUB  x30, x0, x11   // x30 ? 0 - x11 (temp)
    data[14]  = 32'b0111_011110_000000_001011_0000000000;

    // BRN  x6             // if N=1 (ctr>0) loop back
    data[15] = 32'b1011_000000_000110_000000_0000000000;

    // ADD  x10, x0, x5    // result (min) ? x10
    data[18] = 32'b0100_001010_000000_000101_0000000000;
 
    // J    x1             // return to x1
    data[19] = 32'b1000_000000_000001_000000_0000000000;
    */
    
    data[0] = 32'b0100_000001_000001_000010_0000000000;

    data[1] = 32'b0110_000001_000001_0000000000000000;
    
    data[4] = 32'b0011_000000_000100_000001_0000000000;
    
    // SVPC x1, 32
    //data[0] = 32'b1111_000001_0000000000000000100000;
    // ADD x0, x0
    //data[2] = 32'b0111_000000_000000_000000_0000000000;
    // BRZ x1
    //data[3] = 32'b1001_000000_000001_000000_0000000000;
    //data[3] = 32'b1000_000000_000001_0000000000000000;
    //data[3] = 32'b1010_000000_000001_000000_0000000000;
end
assign OUT = data[Address];
endmodule